* SPICE3 file created from NOT_magic.ext - technology: scmos

.option scale=0.09u

M1000 out in VDD w_0_0# pfet w=8 l=2
+  ad=40 pd=26 as=40 ps=26
M1001 out in GND Gnd nfet w=4 l=2
+  ad=20 pd=18 as=29 ps=22
C0 out in 0.05fF
C1 GND in 0.07fF
C2 VDD w_0_0# 0.05fF
C3 out w_0_0# 0.03fF
C4 out VDD 0.11fF
C5 in w_0_0# 0.06fF
C6 VDD in 0.02fF
C7 out GND 0.04fF
C8 GND Gnd 0.16fF
C9 out Gnd 0.05fF
C10 VDD Gnd 0.06fF
C11 in Gnd 0.13fF
C12 w_0_0# Gnd 0.48fF
