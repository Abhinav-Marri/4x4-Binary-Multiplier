magic
tech scmos
timestamp 1669670940
<< polysilicon >>
rect 18 50 62 52
rect 18 26 20 50
rect 26 -55 28 -12
rect 69 -55 71 -51
rect 26 -57 71 -55
<< metal1 >>
rect 13 67 49 71
rect 81 67 124 71
rect 13 35 16 67
rect 120 35 124 67
rect 60 10 64 24
rect 0 6 7 10
rect 38 6 64 10
rect 78 10 81 24
rect 78 6 92 10
rect 124 6 128 10
rect 0 -12 18 -8
rect 47 -8 53 -4
rect 36 -29 39 -12
rect 103 -29 107 -12
rect 36 -33 50 -29
rect 82 -32 107 -29
<< m2contact >>
rect 39 31 45 37
rect 42 -9 47 -4
<< metal2 >>
rect 7 -36 12 -2
rect 42 -4 45 31
rect 49 30 54 34
rect 49 27 57 30
rect 52 3 57 27
rect 52 -2 92 3
rect 7 -41 50 -36
rect 7 -58 12 -41
rect 92 -58 97 -2
rect 7 -63 97 -58
use NAND_magic  NAND_magic_3
timestamp 1669662301
transform 1 0 50 0 1 -28
box 0 -24 32 24
use NAND_magic  NAND_magic_2
timestamp 1669662301
transform 1 0 92 0 1 11
box 0 -24 32 24
use NAND_magic  NAND_magic_1
timestamp 1669662301
transform 1 0 49 0 1 47
box 0 -24 32 24
use NAND_magic  NAND_magic_0
timestamp 1669662301
transform 1 0 7 0 1 11
box 0 -24 32 24
<< labels >>
rlabel metal1 3 8 3 8 3 A
rlabel metal1 3 -10 3 -10 3 B
rlabel metal1 126 8 126 8 7 out
<< end >>
