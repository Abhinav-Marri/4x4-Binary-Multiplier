* SPICE3 file created from OR_magic.ext - technology: scmos

.option scale=0.09u

M1000 NOT_magic_0/in B NOR_magic_0/a_13_6# NOT_magic_0/w_0_0# pfet w=8 l=2
+  ad=40 pd=26 as=48 ps=28
M1001 NOR_magic_0/a_13_6# A VDD NOT_magic_0/w_0_0# pfet w=8 l=2
+  ad=0 pd=0 as=80 ps=52
M1002 GND B NOT_magic_0/in Gnd nfet w=4 l=2
+  ad=87 pd=66 as=24 ps=20
M1003 NOT_magic_0/in A GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 out NOT_magic_0/in VDD NOT_magic_0/w_0_0# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1005 out NOT_magic_0/in GND Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
C0 NOT_magic_0/in VDD 0.10fF
C1 B NOT_magic_0/w_0_0# 0.06fF
C2 GND A 0.07fF
C3 B NOT_magic_0/in 0.10fF
C4 A VDD 0.02fF
C5 NOT_magic_0/in NOT_magic_0/w_0_0# 0.10fF
C6 GND out 0.04fF
C7 B A 0.08fF
C8 out VDD 0.11fF
C9 A NOT_magic_0/w_0_0# 0.06fF
C10 GND B 0.13fF
C11 NOT_magic_0/in A 0.05fF
C12 out NOT_magic_0/w_0_0# 0.03fF
C13 GND NOT_magic_0/in 0.22fF
C14 VDD NOT_magic_0/w_0_0# 0.11fF
C15 out NOT_magic_0/in 0.05fF
C16 out Gnd 0.07fF
C17 GND Gnd 0.38fF
C18 NOT_magic_0/in Gnd 0.20fF
C19 VDD Gnd 0.14fF
C20 B Gnd 0.23fF
C21 A Gnd 0.16fF
C22 NOT_magic_0/w_0_0# Gnd 1.12fF
