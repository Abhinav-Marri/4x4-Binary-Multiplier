* SPICE3 file created from NAND_magic.ext - technology: scmos

.option scale=0.09u

M1000 VDD B out w_0_0# pfet w=8 l=2
+  ad=80 pd=52 as=48 ps=28
M1001 out A VDD w_0_0# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 out B a_13_n12# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1003 a_13_n12# A GND Gnd nfet w=4 l=2
+  ad=0 pd=0 as=29 ps=22
C0 A GND 0.07fF
C1 out w_0_0# 0.02fF
C2 A VDD 0.02fF
C3 A out 0.05fF
C4 B out 0.08fF
C5 VDD out 0.22fF
C6 A w_0_0# 0.06fF
C7 B w_0_0# 0.06fF
C8 VDD w_0_0# 0.09fF
C9 A B 0.08fF
