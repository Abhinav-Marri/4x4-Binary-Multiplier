magic
tech scmos
timestamp 1669709031
<< metal1 >>
rect -83 25 1 29
rect 68 25 73 29
rect -77 -763 -73 -576
rect -69 -617 -65 -364
rect -61 -505 -57 -318
rect -53 -423 -49 -170
rect -45 -229 -41 -106
rect -77 -893 -73 -768
rect -69 -811 -65 -622
rect -61 -699 -57 -510
rect -53 -681 -49 -428
rect -45 -487 -41 -234
rect -37 -247 -33 -60
rect -29 -119 -25 6
rect -29 -183 -25 -124
rect -37 -441 -33 -252
rect -29 -377 -25 -188
rect -22 -37 -18 25
rect -10 7 0 11
rect 70 -16 107 -12
rect -22 -41 2 -37
rect 68 -41 96 -37
rect -22 -295 -18 -41
rect -10 -59 2 -55
rect 300 -73 305 -68
rect 88 -101 93 -95
rect -10 -105 2 -101
rect 68 -105 93 -101
rect 46 -116 50 -113
rect -10 -123 2 -119
rect 46 -120 135 -116
rect 603 -132 607 -12
rect 70 -144 398 -140
rect 871 -151 1390 -145
rect -10 -169 2 -165
rect 68 -169 387 -165
rect -10 -187 2 -183
rect 70 -208 110 -204
rect -10 -233 2 -229
rect 68 -233 99 -229
rect -10 -251 2 -247
rect 366 -265 371 -205
rect 308 -269 371 -265
rect 993 -271 1216 -270
rect 881 -274 1216 -271
rect 993 -275 1216 -274
rect 1384 -280 1390 -151
rect 1481 -282 1619 -280
rect 91 -295 96 -283
rect 1481 -285 1626 -282
rect -22 -299 2 -295
rect 68 -299 96 -295
rect -77 -957 -73 -898
rect -69 -939 -65 -816
rect -61 -829 -57 -704
rect -53 -875 -49 -686
rect -45 -745 -41 -492
rect -37 -635 -33 -446
rect -22 -553 -18 -299
rect -10 -317 1 -313
rect 46 -317 51 -307
rect 46 -322 139 -317
rect 340 -319 975 -313
rect 70 -338 403 -333
rect -10 -363 2 -359
rect 68 -363 258 -359
rect 398 -363 403 -338
rect 969 -344 975 -319
rect 969 -350 981 -344
rect 603 -351 607 -350
rect -10 -381 2 -377
rect 253 -384 258 -363
rect 253 -388 387 -384
rect 1491 -413 1543 -410
rect -10 -427 2 -423
rect 68 -427 332 -422
rect -10 -445 1 -441
rect 70 -466 117 -462
rect -10 -491 2 -487
rect 68 -491 106 -487
rect -10 -509 2 -505
rect 382 -522 387 -442
rect 874 -493 1217 -489
rect 314 -527 387 -522
rect 98 -553 103 -545
rect -22 -557 2 -553
rect 68 -557 103 -553
rect 46 -570 50 -565
rect -10 -575 2 -571
rect 46 -575 145 -570
rect 1213 -572 1217 -493
rect 1540 -506 1543 -413
rect 1619 -441 1626 -285
rect 1787 -504 1792 -500
rect 1540 -510 1570 -506
rect 373 -585 409 -580
rect 882 -584 1008 -581
rect 373 -591 379 -585
rect 70 -596 379 -591
rect 361 -610 398 -605
rect 361 -616 366 -610
rect -10 -621 2 -617
rect 68 -621 366 -616
rect -10 -639 2 -635
rect 390 -681 395 -662
rect 1481 -675 1613 -668
rect -10 -685 2 -681
rect 68 -685 395 -681
rect -10 -703 2 -699
rect 1519 -711 1525 -710
rect 1491 -714 1525 -711
rect -10 -749 2 -745
rect 68 -749 871 -745
rect -10 -767 2 -763
rect 888 -778 892 -715
rect 617 -783 892 -778
rect 70 -790 419 -786
rect 412 -791 419 -790
rect -11 -815 2 -811
rect 68 -815 406 -810
rect -11 -833 2 -829
rect 1519 -844 1525 -714
rect 1607 -781 1613 -675
rect 1782 -771 1787 -674
rect 1519 -849 1550 -844
rect -11 -879 2 -875
rect 68 -879 398 -874
rect 884 -880 1041 -874
rect -11 -897 2 -893
rect 895 -925 1004 -922
rect -11 -943 2 -939
rect 68 -943 421 -936
rect -77 -961 2 -957
rect 415 -1030 421 -943
rect 999 -989 1004 -925
rect 1034 -966 1041 -880
rect 2060 -913 2066 -909
rect 1215 -957 1506 -954
rect 1498 -959 1506 -957
rect 2061 -959 2066 -913
rect 1498 -966 2066 -959
rect 415 -1035 983 -1030
rect 1493 -1100 1500 -1095
<< m2contact >>
rect 65 50 70 55
rect -30 6 -25 11
rect -38 -60 -33 -55
rect -46 -106 -41 -101
rect -54 -170 -49 -165
rect -62 -318 -57 -313
rect -70 -364 -65 -359
rect -78 -576 -73 -571
rect -46 -234 -41 -229
rect -54 -428 -49 -423
rect -62 -510 -57 -505
rect -70 -622 -65 -617
rect -78 -768 -73 -763
rect -30 -124 -25 -119
rect -30 -188 -25 -183
rect -38 -252 -33 -247
rect -30 -382 -25 -377
rect -15 6 -10 11
rect 65 -16 70 -11
rect 602 -12 607 -7
rect -15 -60 -10 -55
rect 65 -80 70 -75
rect -15 -106 -10 -101
rect -15 -124 -10 -119
rect 135 -120 141 -114
rect 65 -144 70 -139
rect -15 -170 -10 -165
rect -15 -188 -10 -183
rect 65 -208 70 -203
rect -15 -234 -10 -229
rect -15 -252 -10 -247
rect 65 -274 70 -269
rect -38 -446 -33 -441
rect -46 -492 -41 -487
rect -54 -686 -49 -681
rect -62 -704 -57 -699
rect -70 -816 -65 -811
rect -78 -898 -73 -893
rect -62 -834 -57 -829
rect -15 -318 -10 -313
rect 139 -322 144 -317
rect 333 -320 340 -313
rect 65 -338 70 -333
rect -15 -364 -10 -359
rect 602 -350 609 -344
rect -15 -382 -10 -377
rect 65 -402 70 -397
rect -15 -428 -10 -423
rect 332 -427 339 -420
rect -15 -446 -10 -441
rect 65 -466 70 -461
rect -15 -492 -10 -487
rect -15 -510 -10 -505
rect 65 -532 70 -527
rect -15 -576 -10 -571
rect 145 -575 151 -569
rect 613 -574 618 -568
rect 65 -596 70 -591
rect -15 -622 -10 -617
rect -38 -640 -33 -635
rect -15 -640 -10 -635
rect 976 -650 981 -645
rect 65 -660 70 -655
rect -15 -686 -10 -681
rect -15 -704 -10 -699
rect 65 -724 70 -719
rect -46 -750 -41 -745
rect -15 -750 -10 -745
rect 871 -749 876 -744
rect -15 -768 -10 -763
rect 65 -790 70 -785
rect -16 -816 -11 -811
rect -16 -834 -11 -829
rect 1782 -674 1787 -667
rect 65 -854 70 -849
rect -54 -880 -49 -875
rect -16 -880 -11 -875
rect -16 -898 -11 -893
rect 65 -918 70 -913
rect -70 -944 -65 -939
rect -16 -944 -11 -939
<< metal2 >>
rect -6 17 3 22
rect -83 7 -30 11
rect -25 7 -15 11
rect -6 -44 -1 17
rect -6 -49 3 -44
rect -83 -59 -38 -55
rect -33 -59 -15 -55
rect -83 -105 -46 -101
rect -41 -105 -15 -101
rect -6 -108 -1 -49
rect -6 -113 3 -108
rect -25 -123 -15 -119
rect -83 -169 -54 -165
rect -49 -169 -15 -165
rect -6 -172 -1 -113
rect -6 -177 3 -172
rect -25 -187 -15 -183
rect -41 -233 -15 -229
rect -6 -236 -1 -177
rect -6 -241 3 -236
rect -33 -251 -15 -247
rect -6 -302 -1 -241
rect -6 -307 3 -302
rect -83 -317 -62 -313
rect -57 -317 -15 -313
rect -83 -363 -70 -359
rect -65 -363 -15 -359
rect -6 -366 -1 -307
rect -6 -371 3 -366
rect -25 -381 -15 -377
rect -49 -427 -15 -423
rect -6 -430 -1 -371
rect -6 -435 3 -430
rect -33 -445 -15 -441
rect -41 -491 -15 -487
rect -6 -494 -1 -435
rect -6 -499 3 -494
rect -57 -509 -15 -505
rect -6 -560 -1 -499
rect -6 -565 3 -560
rect -83 -575 -78 -571
rect -73 -575 -15 -571
rect -65 -621 -15 -617
rect -6 -624 -1 -565
rect -6 -629 3 -624
rect -33 -639 -15 -635
rect -49 -685 -15 -681
rect -6 -688 -1 -629
rect -6 -693 3 -688
rect -57 -703 -15 -699
rect -41 -749 -15 -745
rect -6 -752 -1 -693
rect -6 -757 3 -752
rect -73 -767 -15 -763
rect -65 -815 -16 -811
rect -6 -818 -1 -757
rect -6 -823 3 -818
rect -57 -833 -16 -829
rect -49 -879 -16 -875
rect -6 -882 -1 -823
rect -6 -887 3 -882
rect -73 -897 -16 -893
rect -65 -943 -16 -939
rect -6 -946 -1 -887
rect 70 -918 74 54
rect 173 -10 602 -7
rect 265 -181 270 -146
rect 265 -186 366 -181
rect 175 -203 356 -199
rect 268 -432 273 -338
rect 333 -420 339 -320
rect 351 -345 356 -203
rect 362 -229 366 -186
rect 884 -205 889 -200
rect 362 -235 434 -229
rect 1494 -344 1499 -339
rect 351 -350 602 -345
rect 997 -419 1002 -344
rect 884 -424 1002 -419
rect 268 -436 436 -432
rect 183 -455 406 -454
rect 183 -457 407 -455
rect 183 -459 187 -457
rect 402 -537 407 -457
rect 1046 -502 1052 -412
rect 1655 -434 1803 -430
rect 1798 -460 1803 -434
rect 1046 -509 1051 -502
rect 847 -515 1051 -509
rect 402 -542 618 -537
rect 614 -568 618 -542
rect 275 -696 280 -596
rect 895 -618 981 -613
rect 895 -646 901 -618
rect 1578 -639 1583 -504
rect 1493 -645 1585 -639
rect 960 -650 976 -645
rect 275 -703 444 -696
rect 333 -888 339 -703
rect 793 -755 801 -748
rect 960 -745 967 -650
rect 876 -749 967 -745
rect 1041 -755 1047 -713
rect 1632 -741 1642 -573
rect 1798 -668 1802 -460
rect 1787 -673 1803 -668
rect 1798 -676 1802 -673
rect 1437 -749 1642 -741
rect 793 -760 1047 -755
rect 1041 -761 1047 -760
rect 1402 -813 1411 -812
rect 1402 -821 1550 -813
rect 1402 -849 1411 -821
rect 2063 -844 2069 -839
rect 898 -856 1411 -849
rect 333 -894 450 -888
rect -6 -951 3 -946
rect 812 -1067 820 -959
rect 1496 -1030 1503 -1025
rect 812 -1073 1045 -1067
rect 1611 -1117 1618 -913
rect 1459 -1123 1618 -1117
use AND_magic  AND_magic_15
timestamp 1669670829
transform 1 0 3 0 1 -957
box -3 -11 65 43
use FA_magic  FA_magic_3
timestamp 1669671046
transform 1 0 432 0 1 -975
box -47 16 466 192
use AND_magic  AND_magic_14
timestamp 1669670829
transform 1 0 3 0 1 -893
box -3 -11 65 43
use FA_magic  FA_magic_4
timestamp 1669671046
transform 1 0 1030 0 1 -1149
box -47 16 466 192
use FA_magic  FA_magic_7
timestamp 1669671046
transform 1 0 1597 0 1 -963
box -47 16 466 192
use AND_magic  AND_magic_13
timestamp 1669670829
transform 1 0 3 0 1 -829
box -3 -11 65 43
use AND_magic  AND_magic_12
timestamp 1669670829
transform 1 0 3 0 1 -763
box -3 -11 65 43
use AND_magic  AND_magic_11
timestamp 1669670829
transform 1 0 3 0 1 -699
box -3 -11 65 43
use FA_magic  FA_magic_2
timestamp 1669671046
transform 1 0 429 0 1 -765
box -47 16 466 192
use FA_magic  FA_magic_6
timestamp 1669671046
transform 1 0 1028 0 1 -764
box -47 16 466 192
use AND_magic  AND_magic_10
timestamp 1669670829
transform 1 0 3 0 1 -635
box -3 -11 65 43
use HA_magic  HA_magic_2
timestamp 1669670993
transform 1 0 61 0 1 -586
box 37 -10 254 129
use AND_magic  AND_magic_9
timestamp 1669670829
transform 1 0 3 0 1 -571
box -3 -11 65 43
use AND_magic  AND_magic_8
timestamp 1669670829
transform 1 0 3 0 1 -505
box -3 -11 65 43
use AND_magic  AND_magic_7
timestamp 1669670829
transform 1 0 3 0 1 -441
box -3 -11 65 43
use FA_magic  FA_magic_1
timestamp 1669671046
transform 1 0 418 0 1 -543
box -47 16 466 192
use FA_magic  FA_magic_5
timestamp 1669671046
transform 1 0 1028 0 1 -463
box -47 16 466 192
use HA_magic  HA_magic_3
timestamp 1669670993
transform 1 0 1533 0 1 -563
box 37 -10 254 129
use AND_magic  AND_magic_6
timestamp 1669670829
transform 1 0 3 0 1 -377
box -3 -11 65 43
use HA_magic  HA_magic_1
timestamp 1669670993
transform 1 0 54 0 1 -328
box 37 -10 254 129
use AND_magic  AND_magic_5
timestamp 1669670829
transform 1 0 3 0 1 -313
box -3 -11 65 43
use AND_magic  AND_magic_4
timestamp 1669670829
transform 1 0 3 0 1 -247
box -3 -11 65 43
use FA_magic  FA_magic_0
timestamp 1669671046
transform 1 0 418 0 1 -324
box -47 16 466 192
use AND_magic  AND_magic_3
timestamp 1669670829
transform 1 0 3 0 1 -183
box -3 -11 65 43
use HA_magic  HA_magic_0
timestamp 1669670993
transform 1 0 51 0 1 -136
box 37 -10 254 129
use AND_magic  AND_magic_2
timestamp 1669670829
transform 1 0 3 0 1 -119
box -3 -11 65 43
use AND_magic  AND_magic_1
timestamp 1669670829
transform 1 0 3 0 1 -55
box -3 -11 65 43
use AND_magic  AND_magic_0
timestamp 1669670829
transform 1 0 3 0 1 11
box -3 -11 65 43
<< labels >>
rlabel metal2 -83 -575 -79 -571 3 B3
rlabel metal2 -83 -363 -79 -359 3 A3
rlabel metal2 -83 -317 -79 -313 3 B2
rlabel metal2 -83 -169 -79 -165 3 A2
rlabel metal2 -83 -105 -79 -101 3 A1
rlabel metal2 -83 -59 -79 -55 3 B1
rlabel metal1 -83 25 -79 29 3 A0
rlabel metal2 -83 7 -79 11 3 B0
rlabel metal1 68 25 73 29 7 P0
rlabel metal1 300 -73 305 -68 7 P1
rlabel metal2 884 -205 889 -200 7 P2
rlabel metal2 1494 -344 1499 -339 7 P3
rlabel metal1 1787 -504 1792 -500 7 P4
rlabel metal2 2063 -844 2069 -839 7 P5
rlabel metal2 1496 -1030 1503 -1025 1 P6
rlabel metal1 1493 -1100 1500 -1095 1 C5
<< end >>
