magic
tech scmos
timestamp 1669662021
<< nwell >>
rect 0 0 24 20
<< ntransistor >>
rect 11 -12 13 -8
<< ptransistor >>
rect 11 6 13 14
<< ndiffusion >>
rect 10 -12 11 -8
rect 13 -12 14 -8
<< pdiffusion >>
rect 10 6 11 14
rect 13 6 14 14
<< ndcontact >>
rect 14 -12 18 -8
<< pdcontact >>
rect 6 6 10 14
rect 14 6 18 14
<< polysilicon >>
rect 11 14 13 17
rect 11 -8 13 6
rect 11 -15 13 -12
<< polycontact >>
rect 7 -5 11 -1
<< metal1 >>
rect 0 20 24 24
rect 6 14 10 20
rect 14 -1 18 6
rect 0 -5 7 -1
rect 14 -5 24 -1
rect 14 -8 18 -5
<< ndm12contact >>
rect 5 -13 10 -8
<< metal2 >>
rect 0 -13 5 -8
<< labels >>
rlabel metal1 0 20 24 24 5 VDD
rlabel metal2 0 -13 5 -8 2 GND
rlabel metal1 21 -3 21 -3 7 out
rlabel metal1 3 -3 3 -3 3 in
<< end >>
